`ifndef PERIOD
`define PERIOD 10
`endif

`ifndef CYCLES
`define CYCLES 1000000
`endif

`ifndef OUTPUT
`define OUTPUT "audio_output_test.vcd"
`endif
