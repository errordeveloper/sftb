module main;

initial $sftb_open_input_file;

initial begin
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
#10 $sftb_fetch_sample();
end

endmodule
