module main;

initial $sftb_open_input_file;

initial $sftb_fetch_sample;

endmodule
